`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:32:32 04/02/2018 
// Design Name: 
// Module Name:    ksablocking1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ksablocking1(
    input reset,
    input write_en,
    input clock,
    input [31:0] fp_input,
    input [7:0] input_length,
    output [31:0] sum
    );

	
	
	
endmodule
